module vpcie_header (
        output reg [7:0] op
    );
endmodule // vpcie_header
